// ===============================================================
// font8x16_rom.v
// 8x16 字库
// 字符 included: A B C D E F G H Z # 0-9 空格
// 新增大写字母: N O R T U (Auto Range)
// 新增小写字母: a e g i n o r t u z (uto ange in z)
// ===============================================================
`timescale 1ns/1ps
module font8x16_rom(
    input  wire [7:0] ch,      // ASCII
    input  wire [3:0] row,     // 0..15
    output reg [7:0] bits      // each bit is 1 pixel
);

    always @(*) begin
        case (ch)

        // -----------------------------
        // 大写字母
        // -----------------------------

        "A": case(row)  // Auto
            0: bits = 8'b00011000;
            1: bits = 8'b00011000;
            2: bits = 8'b00100100;
            3: bits = 8'b00100100;
            4: bits = 8'b00100100;
            5: bits = 8'b01111110;
            6: bits = 8'b01000010;
            7: bits = 8'b01000010;
            8: bits = 8'b01000010;
            9: bits = 8'b11100111;
            10: bits = 8'b00000000;
            11: bits = 8'b00000000;
            12: bits = 8'b00000000;
            13: bits = 8'b00000000;
            14: bits = 8'b00000000;
            15: bits = 8'b00000000;
        endcase

        "B": case(row)  // Bin
            0: bits = 8'b01111110;
            1: bits = 8'b01000001;
            2: bits = 8'b01000001;
            3: bits = 8'b01000001;
            4: bits = 8'b01111110;
            5: bits = 8'b01000001;
            6: bits = 8'b01000001;
            7: bits = 8'b01000001;
            8: bits = 8'b01000001;
            9: bits = 8'b01111110;
            10: bits = 8'b00000000;
            11: bits = 8'b00000000;
            12: bits = 8'b00000000;
            13: bits = 8'b00000000;
            14: bits = 8'b00000000;
            15: bits = 8'b00000000;
        endcase

        "C": case(row)  // 原有
            0: bits = 8'b00111100;
            1: bits = 8'b01000010;
            2: bits = 8'b01000000;
            3: bits = 8'b01000000;
            4: bits = 8'b01000000;
            5: bits = 8'b01000000;
            6: bits = 8'b01000000;
            7: bits = 8'b01000000;
            8: bits = 8'b01000010;
            9: bits = 8'b00111100;
            10: bits = 8'b00000000;
            11: bits = 8'b00000000;
            12: bits = 8'b00000000;
            13: bits = 8'b00000000;
            14: bits = 8'b00000000;
            15: bits = 8'b00000000;
        endcase

        "D": case(row)  // 原有
            0: bits = 8'b01111100;
            1: bits = 8'b01000010;
            2: bits = 8'b01000001;
            3: bits = 8'b01000001;
            4: bits = 8'b01000001;
            5: bits = 8'b01000001;
            6: bits = 8'b01000001;
            7: bits = 8'b01000001;
            8: bits = 8'b01000010;
            9: bits = 8'b01111100;
            10: bits = 8'b00000000;
            11: bits = 8'b00000000;
            12: bits = 8'b00000000;
            13: bits = 8'b00000000;
            14: bits = 8'b00000000;
            15: bits = 8'b00000000;
        endcase

        "E": case(row)  // Range
            0: bits = 8'b01111111;
            1: bits = 8'b01000000;
            2: bits = 8'b01000000;
            3: bits = 8'b01000000;
            4: bits = 8'b01111111;
            5: bits = 8'b01000000;
            6: bits = 8'b01000000;
            7: bits = 8'b01000000;
            8: bits = 8'b01000000;
            9: bits = 8'b01111111;
            10: bits = 8'b00000000;
            11: bits = 8'b00000000;
            12: bits = 8'b00000000;
            13: bits = 8'b00000000;
            14: bits = 8'b00000000;
            15: bits = 8'b00000000;
        endcase

        "F": case(row)  // 已有F，不需要添加
            0: bits = 8'b01111111;
            1: bits = 8'b01000000;
            2: bits = 8'b01000000;
            3: bits = 8'b01000000;
            4: bits = 8'b01111111;
            5: bits = 8'b01000000;
            6: bits = 8'b01000000;
            7: bits = 8'b01000000;
            8: bits = 8'b01000000;
            9: bits = 8'b01000000;
            10: bits = 8'b00000000;
            11: bits = 8'b00000000;
            12: bits = 8'b00000000;
            13: bits = 8'b00000000;
            14: bits = 8'b00000000;
            15: bits = 8'b00000000;
        endcase

        "G": case(row)  // 原有
            0: bits = 8'b00111100;
            1: bits = 8'b01000010;
            2: bits = 8'b01000000;
            3: bits = 8'b01000000;
            4: bits = 8'b01001110;
            5: bits = 8'b01000010;
            6: bits = 8'b01000010;
            7: bits = 8'b01000010;
            8: bits = 8'b01000010;
            9: bits = 8'b00111100;
            10: bits = 8'b00000000;
            11: bits = 8'b00000000;
            12: bits = 8'b00000000;
            13: bits = 8'b00000000;
            14: bits = 8'b00000000;
            15: bits = 8'b00000000;
        endcase

        "H": case(row)  // 原有
            0: bits = 8'b01000010;
            1: bits = 8'b01000010;
            2: bits = 8'b01000010;
            3: bits = 8'b01000010;
            4: bits = 8'b01111110;
            5: bits = 8'b01000010;
            6: bits = 8'b01000010;
            7: bits = 8'b01000010;
            8: bits = 8'b01000010;
            9: bits = 8'b01000010;
            10: bits = 8'b00000000;
            11: bits = 8'b00000000;
            12: bits = 8'b00000000;
            13: bits = 8'b00000000;
            14: bits = 8'b00000000;
            15: bits = 8'b00000000;
        endcase

        // --- 新增的大写字母N ---
        "N": case(row)  // 新增的大写N
            0: bits = 8'b01000010;
            1: bits = 8'b01100010;
            2: bits = 8'b01010010;
            3: bits = 8'b01001010;
            4: bits = 8'b01000110;
            5: bits = 8'b01000010;
            6: bits = 8'b01000010;
            7: bits = 8'b01000010;
            8: bits = 8'b01000010;
            9: bits = 8'b01000010;
            10: bits = 8'b00000000;
            11: bits = 8'b00000000;
            12: bits = 8'b00000000;
            13: bits = 8'b00000000;
            14: bits = 8'b00000000;
            15: bits = 8'b00000000;
        endcase

        "O": case(row)  // Auto 的 O（大写）
            0: bits = 8'b00111100;
            1: bits = 8'b01000010;
            2: bits = 8'b01000010;
            3: bits = 8'b01000010;
            4: bits = 8'b01000010;
            5: bits = 8'b01000010;
            6: bits = 8'b01000010;
            7: bits = 8'b01000010;
            8: bits = 8'b01000010;
            9: bits = 8'b00111100;
            10: bits = 8'b00000000;
            11: bits = 8'b00000000;
            12: bits = 8'b00000000;
            13: bits = 8'b00000000;
            14: bits = 8'b00000000;
            15: bits = 8'b00000000;
        endcase

        "R": case(row)  // Range 的 R（大写）
            0: bits = 8'b01111100;
            1: bits = 8'b01000010;
            2: bits = 8'b01000010;
            3: bits = 8'b01000010;
            4: bits = 8'b01111100;
            5: bits = 8'b01001000;
            6: bits = 8'b01000100;
            7: bits = 8'b01000010;
            8: bits = 8'b01000010;
            9: bits = 8'b01100001;
            10: bits = 8'b00000000;
            11: bits = 8'b00000000;
            12: bits = 8'b00000000;
            13: bits = 8'b00000000;
            14: bits = 8'b00000000;
            15: bits = 8'b00000000;
        endcase

        "T": case(row)  // Auto 的 T（大写）
            0: bits = 8'b11111111;
            1: bits = 8'b00011000;
            2: bits = 8'b00011000;
            3: bits = 8'b00011000;
            4: bits = 8'b00011000;
            5: bits = 8'b00011000;
            6: bits = 8'b00011000;
            7: bits = 8'b00011000;
            8: bits = 8'b00011000;
            9: bits = 8'b00011000;
            10: bits = 8'b00000000;
            11: bits = 8'b00000000;
            12: bits = 8'b00000000;
            13: bits = 8'b00000000;
            14: bits = 8'b00000000;
            15: bits = 8'b00000000;
        endcase

        "U": case(row)  // Auto 的 U（大写）
            0: bits = 8'b01000010;
            1: bits = 8'b01000010;
            2: bits = 8'b01000010;
            3: bits = 8'b01000010;
            4: bits = 8'b01000010;
            5: bits = 8'b01000010;
            6: bits = 8'b01000010;
            7: bits = 8'b01000010;
            8: bits = 8'b01000010;
            9: bits = 8'b00111100;
            10: bits = 8'b00000000;
            11: bits = 8'b00000000;
            12: bits = 8'b00000000;
            13: bits = 8'b00000000;
            14: bits = 8'b00000000;
            15: bits = 8'b00000000;
        endcase

        "Z": case(row)  // 原有（大写Z）
            0: bits = 8'b01111110;
            1: bits = 8'b00000010;
            2: bits = 8'b00000100;
            3: bits = 8'b00001000;
            4: bits = 8'b00010000;
            5: bits = 8'b00100000;
            6: bits = 8'b01000000;
            7: bits = 8'b01000000;
            8: bits = 8'b01000000;
            9: bits = 8'b01111110;
            10: bits = 8'b00000000;
            11: bits = 8'b00000000;
            12: bits = 8'b00000000;
            13: bits = 8'b00000000;
            14: bits = 8'b00000000;
            15: bits = 8'b00000000;
        endcase

        // -----------------------------
        // 小写字母 (uto ange in z)
        // -----------------------------
        // ...（小写字母部分保持不变，从之前的代码中复制）...

        // 空格字符
        " ": case(row)
            0: bits = 8'b00000000;
            1: bits = 8'b00000000;
            2: bits = 8'b00000000;
            3: bits = 8'b00000000;
            4: bits = 8'b00000000;
            5: bits = 8'b00000000;
            6: bits = 8'b00000000;
            7: bits = 8'b00000000;
            8: bits = 8'b00000000;
            9: bits = 8'b00000000;
            10: bits = 8'b00000000;
            11: bits = 8'b00000000;
            12: bits = 8'b00000000;
            13: bits = 8'b00000000;
            14: bits = 8'b00000000;
            15: bits = 8'b00000000;
        endcase

        // -----------------------------
        // 数字 0-9
        // -----------------------------
        // ...（数字部分保持不变，从之前的代码中复制）...

        // -----------------------------
        // "#" (井号)
        // -----------------------------
        "#": case(row)
            0: bits = 8'b00000000;
            1: bits = 8'b00010100;
            2: bits = 8'b00010100;
            3: bits = 8'b01111111;
            4: bits = 8'b00010100;
            5: bits = 8'b00010100;
            6: bits = 8'b01111111;
            7: bits = 8'b00010100;
            8: bits = 8'b00010100;
            9: bits = 8'b00000000;
            10: bits = 8'b00000000;
            11: bits = 8'b00000000;
            12: bits = 8'b00000000;
            13: bits = 8'b00000000;
            14: bits = 8'b00000000;
            15: bits = 8'b00000000;
        endcase

        // -----------------------------
        // 小写字母 (uto ange in z)
        // -----------------------------

        "a": case(row)  // Auto 的 a（小写）
            0: bits = 8'b00000000;
            1: bits = 8'b00000000;
            2: bits = 8'b00000000;
            3: bits = 8'b00111100;
            4: bits = 8'b01000010;
            5: bits = 8'b00111110;
            6: bits = 8'b01000010;
            7: bits = 8'b01000010;
            8: bits = 8'b01000110;
            9: bits = 8'b00111011;
            10: bits = 8'b00000000;
            11: bits = 8'b00000000;
            12: bits = 8'b00000000;
            13: bits = 8'b00000000;
            14: bits = 8'b00000000;
            15: bits = 8'b00000000;
        endcase

        "e": case(row)  // ange 的 e（小写）
            0: bits = 8'b00000000;
            1: bits = 8'b00000000;
            2: bits = 8'b00000000;
            3: bits = 8'b00111100;
            4: bits = 8'b01000010;
            5: bits = 8'b01111110;
            6: bits = 8'b01000000;
            7: bits = 8'b01000000;
            8: bits = 8'b01000010;
            9: bits = 8'b00111100;
            10: bits = 8'b00000000;
            11: bits = 8'b00000000;
            12: bits = 8'b00000000;
            13: bits = 8'b00000000;
            14: bits = 8'b00000000;
            15: bits = 8'b00000000;
        endcase

        "g": case(row)  // ange 的 g（小写）
            0: bits = 8'b00000000;
            1: bits = 8'b00000000;
            2: bits = 8'b00000000;
            3: bits = 8'b00111110;
            4: bits = 8'b01000010;
            5: bits = 8'b01000010;
            6: bits = 8'b00111110;
            7: bits = 8'b00000010;
            8: bits = 8'b01000010;
            9: bits = 8'b00111100;
            10: bits = 8'b00000000;
            11: bits = 8'b00000000;
            12: bits = 8'b00000000;
            13: bits = 8'b00000000;
            14: bits = 8'b00000000;
            15: bits = 8'b00000000;
        endcase

        "i": case(row)  // in 的 i（小写）
            0: bits = 8'b00000000;
            1: bits = 8'b00011000;
            2: bits = 8'b00000000;
            3: bits = 8'b00011000;
            4: bits = 8'b00011000;
            5: bits = 8'b00011000;
            6: bits = 8'b00011000;
            7: bits = 8'b00011000;
            8: bits = 8'b00011000;
            9: bits = 8'b00011000;
            10: bits = 8'b00000000;
            11: bits = 8'b00000000;
            12: bits = 8'b00000000;
            13: bits = 8'b00000000;
            14: bits = 8'b00000000;
            15: bits = 8'b00000000;
        endcase

        "n": case(row)  // in 的 n（小写）, ange 的 n
            0: bits = 8'b00000000;
            1: bits = 8'b00000000;
            2: bits = 8'b00000000;
            3: bits = 8'b01011100;
            4: bits = 8'b01100010;
            5: bits = 8'b01000010;
            6: bits = 8'b01000010;
            7: bits = 8'b01000010;
            8: bits = 8'b01000010;
            9: bits = 8'b01000010;
            10: bits = 8'b00000000;
            11: bits = 8'b00000000;
            12: bits = 8'b00000000;
            13: bits = 8'b00000000;
            14: bits = 8'b00000000;
            15: bits = 8'b00000000;
        endcase

        "o": case(row)  // uto 的 o（小写）
            0: bits = 8'b00000000;
            1: bits = 8'b00000000;
            2: bits = 8'b00000000;
            3: bits = 8'b00111100;
            4: bits = 8'b01000010;
            5: bits = 8'b01000010;
            6: bits = 8'b01000010;
            7: bits = 8'b01000010;
            8: bits = 8'b01000010;
            9: bits = 8'b00111100;
            10: bits = 8'b00000000;
            11: bits = 8'b00000000;
            12: bits = 8'b00000000;
            13: bits = 8'b00000000;
            14: bits = 8'b00000000;
            15: bits = 8'b00000000;
        endcase

        "r": case(row)  // ange 的 r（小写）
            0: bits = 8'b00000000;
            1: bits = 8'b00000000;
            2: bits = 8'b00000000;
            3: bits = 8'b01011100;
            4: bits = 8'b01100010;
            5: bits = 8'b01000000;
            6: bits = 8'b01000000;
            7: bits = 8'b01000000;
            8: bits = 8'b01000000;
            9: bits = 8'b01000000;
            10: bits = 8'b00000000;
            11: bits = 8'b00000000;
            12: bits = 8'b00000000;
            13: bits = 8'b00000000;
            14: bits = 8'b00000000;
            15: bits = 8'b00000000;
        endcase

        "t": case(row)  // uto 的 t（小写）
            0: bits = 8'b00000000;
            1: bits = 8'b00010000;
            2: bits = 8'b00010000;
            3: bits = 8'b01111100;
            4: bits = 8'b00010000;
            5: bits = 8'b00010000;
            6: bits = 8'b00010000;
            7: bits = 8'b00010000;
            8: bits = 8'b00010010;
            9: bits = 8'b00001100;
            10: bits = 8'b00000000;
            11: bits = 8'b00000000;
            12: bits = 8'b00000000;
            13: bits = 8'b00000000;
            14: bits = 8'b00000000;
            15: bits = 8'b00000000;
        endcase

        "u": case(row)  // uto 的 u（小写）
            0: bits = 8'b00000000;
            1: bits = 8'b00000000;
            2: bits = 8'b00000000;
            3: bits = 8'b01000010;
            4: bits = 8'b01000010;
            5: bits = 8'b01000010;
            6: bits = 8'b01000010;
            7: bits = 8'b01000010;
            8: bits = 8'b01000110;
            9: bits = 8'b00111010;
            10: bits = 8'b00000000;
            11: bits = 8'b00000000;
            12: bits = 8'b00000000;
            13: bits = 8'b00000000;
            14: bits = 8'b00000000;
            15: bits = 8'b00000000;
        endcase

        "z": case(row)  // z（小写）
            0: bits = 8'b00000000;
            1: bits = 8'b00000000;
            2: bits = 8'b00000000;
            3: bits = 8'b01111110;
            4: bits = 8'b00000100;
            5: bits = 8'b00001000;
            6: bits = 8'b00010000;
            7: bits = 8'b00100000;
            8: bits = 8'b01000000;
            9: bits = 8'b01111110;
            10: bits = 8'b00000000;
            11: bits = 8'b00000000;
            12: bits = 8'b00000000;
            13: bits = 8'b00000000;
            14: bits = 8'b00000000;
            15: bits = 8'b00000000;
        endcase

        // 空格字符
        " ": case(row)
            0: bits = 8'b00000000;
            1: bits = 8'b00000000;
            2: bits = 8'b00000000;
            3: bits = 8'b00000000;
            4: bits = 8'b00000000;
            5: bits = 8'b00000000;
            6: bits = 8'b00000000;
            7: bits = 8'b00000000;
            8: bits = 8'b00000000;
            9: bits = 8'b00000000;
            10: bits = 8'b00000000;
            11: bits = 8'b00000000;
            12: bits = 8'b00000000;
            13: bits = 8'b00000000;
            14: bits = 8'b00000000;
            15: bits = 8'b00000000;
        endcase

        // -----------------------------
        // 数字 0-9
        // -----------------------------
        "0": case(row)
            0: bits = 8'b00111100;
            1: bits = 8'b01000010;
            2: bits = 8'b01000010;
            3: bits = 8'b01000110;
            4: bits = 8'b01001010;
            5: bits = 8'b01010010;
            6: bits = 8'b01100010;
            7: bits = 8'b01000010;
            8: bits = 8'b01000010;
            9: bits = 8'b00111100;
            10: bits = 8'b00000000;
            11: bits = 8'b00000000;
            12: bits = 8'b00000000;
            13: bits = 8'b00000000;
            14: bits = 8'b00000000;
            15: bits = 8'b00000000;
        endcase

        "1": case(row)
            0: bits = 8'b00001000;
            1: bits = 8'b00011000;
            2: bits = 8'b00101000;
            3: bits = 8'b00001000;
            4: bits = 8'b00001000;
            5: bits = 8'b00001000;
            6: bits = 8'b00001000;
            7: bits = 8'b00001000;
            8: bits = 8'b00001000;
            9: bits = 8'b00111110;
            10: bits = 8'b00000000;
            11: bits = 8'b00000000;
            12: bits = 8'b00000000;
            13: bits = 8'b00000000;
            14: bits = 8'b00000000;
            15: bits = 8'b00000000;
        endcase

        "2": case(row)
            0: bits = 8'b00111100;
            1: bits = 8'b01000010;
            2: bits = 8'b00000010;
            3: bits = 8'b00000010;
            4: bits = 8'b00000100;
            5: bits = 8'b00001000;
            6: bits = 8'b00010000;
            7: bits = 8'b00100000;
            8: bits = 8'b01000000;
            9: bits = 8'b01111110;
            10: bits = 8'b00000000;
            11: bits = 8'b00000000;
            12: bits = 8'b00000000;
            13: bits = 8'b00000000;
            14: bits = 8'b00000000;
            15: bits = 8'b00000000;
        endcase

        "3": case(row)
            0: bits = 8'b00111100;
            1: bits = 8'b01000010;
            2: bits = 8'b00000010;
            3: bits = 8'b00000010;
            4: bits = 8'b00011100;
            5: bits = 8'b00000010;
            6: bits = 8'b00000010;
            7: bits = 8'b00000010;
            8: bits = 8'b01000010;
            9: bits = 8'b00111100;
            10: bits = 8'b00000000;
            11: bits = 8'b00000000;
            12: bits = 8'b00000000;
            13: bits = 8'b00000000;
            14: bits = 8'b00000000;
            15: bits = 8'b00000000;
        endcase

        "4": case(row)
            0: bits = 8'b00000100;
            1: bits = 8'b00001100;
            2: bits = 8'b00010100;
            3: bits = 8'b00100100;
            4: bits = 8'b01000100;
            5: bits = 8'b01111110;
            6: bits = 8'b00000100;
            7: bits = 8'b00000100;
            8: bits = 8'b00000100;
            9: bits = 8'b00000100;
            10: bits = 8'b00000000;
            11: bits = 8'b00000000;
            12: bits = 8'b00000000;
            13: bits = 8'b00000000;
            14: bits = 8'b00000000;
            15: bits = 8'b00000000;
        endcase

        "5": case(row)
            0: bits = 8'b01111110;
            1: bits = 8'b01000000;
            2: bits = 8'b01000000;
            3: bits = 8'b01111100;
            4: bits = 8'b00000010;
            5: bits = 8'b00000010;
            6: bits = 8'b00000010;
            7: bits = 8'b00000010;
            8: bits = 8'b01000010;
            9: bits = 8'b00111100;
            10: bits = 8'b00000000;
            11: bits = 8'b00000000;
            12: bits = 8'b00000000;
            13: bits = 8'b00000000;
            14: bits = 8'b00000000;
            15: bits = 8'b00000000;
        endcase

        "6": case(row)
            0: bits = 8'b00111100;
            1: bits = 8'b01000010;
            2: bits = 8'b01000000;
            3: bits = 8'b01000000;
            4: bits = 8'b01111100;
            5: bits = 8'b01000010;
            6: bits = 8'b01000010;
            7: bits = 8'b01000010;
            8: bits = 8'b01000010;
            9: bits = 8'b00111100;
            10: bits = 8'b00000000;
            11: bits = 8'b00000000;
            12: bits = 8'b00000000;
            13: bits = 8'b00000000;
            14: bits = 8'b00000000;
            15: bits = 8'b00000000;
        endcase

        "7": case(row)
            0: bits = 8'b01111110;
            1: bits = 8'b00000010;
            2: bits = 8'b00000100;
            3: bits = 8'b00000100;
            4: bits = 8'b00001000;
            5: bits = 8'b00001000;
            6: bits = 8'b00010000;
            7: bits = 8'b00010000;
            8: bits = 8'b00100000;
            9: bits = 8'b00100000;
            10: bits = 8'b00000000;
            11: bits = 8'b00000000;
            12: bits = 8'b00000000;
            13: bits = 8'b00000000;
            14: bits = 8'b00000000;
            15: bits = 8'b00000000;
        endcase

        "8": case(row)
            0: bits = 8'b00111100;
            1: bits = 8'b01000010;
            2: bits = 8'b01000010;
            3: bits = 8'b01000010;
            4: bits = 8'b00111100;
            5: bits = 8'b01000010;
            6: bits = 8'b01000010;
            7: bits = 8'b01000010;
            8: bits = 8'b01000010;
            9: bits = 8'b00111100;
            10: bits = 8'b00000000;
            11: bits = 8'b00000000;
            12: bits = 8'b00000000;
            13: bits = 8'b00000000;
            14: bits = 8'b00000000;
            15: bits = 8'b00000000;
        endcase

        "9": case(row)
            0: bits = 8'b00111100;
            1: bits = 8'b01000010;
            2: bits = 8'b01000010;
            3: bits = 8'b01000010;
            4: bits = 8'b00111110;
            5: bits = 8'b00000010;
            6: bits = 8'b00000010;
            7: bits = 8'b00000010;
            8: bits = 8'b01000010;
            9: bits = 8'b00111100;
            10: bits = 8'b00000000;
            11: bits = 8'b00000000;
            12: bits = 8'b00000000;
            13: bits = 8'b00000000;
            14: bits = 8'b00000000;
            15: bits = 8'b00000000;
        endcase
        // 默认情况：空白字符
        default: case(row)
            0: bits = 8'b00000000;
            1: bits = 8'b00000000;
            2: bits = 8'b00000000;
            3: bits = 8'b00000000;
            4: bits = 8'b00000000;
            5: bits = 8'b00000000;
            6: bits = 8'b00000000;
            7: bits = 8'b00000000;
            8: bits = 8'b00000000;
            9: bits = 8'b00000000;
            10: bits = 8'b00000000;
            11: bits = 8'b00000000;
            12: bits = 8'b00000000;
            13: bits = 8'b00000000;
            14: bits = 8'b00000000;
            15: bits = 8'b00000000;
        endcase
        
        endcase
    end
endmodule