
`ifndef HANN_WINDOW_COEFF_SV
`define HANN_WINDOW_COEFF_SV

package hann_window_coeff;
localparam [15:0] HANN_128 [0:127] = '{
    16'h0000, 16'h0014, 16'h0050, 16'h00B4, 16'h013F, 16'h01F2, 16'h02CC, 16'h03CC, 
    16'h04F2, 16'h063D, 16'h07AC, 16'h093E, 16'h0AF3, 16'h0CC9, 16'h0EBF, 16'h10D4, 
    16'h1306, 16'h1555, 16'h17BE, 16'h1A40, 16'h1CDA, 16'h1F8B, 16'h224F, 16'h2526, 
    16'h280E, 16'h2B05, 16'h2E09, 16'h3118, 16'h3431, 16'h3751, 16'h3A76, 16'h3D9F, 
    16'h40CA, 16'h43F4, 16'h471B, 16'h4A3E, 16'h4D5B, 16'h506F, 16'h5379, 16'h5676, 
    16'h5966, 16'h5C46, 16'h5F14, 16'h61CE, 16'h6474, 16'h6702, 16'h6978, 16'h6BD4, 
    16'h6E15, 16'h7039, 16'h723E, 16'h7424, 16'h75EA, 16'h778D, 16'h790E, 16'h7A6B, 
    16'h7BA4, 16'h7CB7, 16'h7DA4, 16'h7E6A, 16'h7F09, 16'h7F81, 16'h7FD1, 16'h7FF9, 
    16'h7FF9, 16'h7FD1, 16'h7F81, 16'h7F09, 16'h7E6A, 16'h7DA4, 16'h7CB7, 16'h7BA4, 
    16'h7A6B, 16'h790E, 16'h778D, 16'h75EA, 16'h7424, 16'h723E, 16'h7039, 16'h6E15, 
    16'h6BD4, 16'h6978, 16'h6702, 16'h6474, 16'h61CE, 16'h5F14, 16'h5C46, 16'h5966, 
    16'h5676, 16'h5379, 16'h506F, 16'h4D5B, 16'h4A3E, 16'h471B, 16'h43F4, 16'h40CA, 
    16'h3D9F, 16'h3A76, 16'h3751, 16'h3431, 16'h3118, 16'h2E09, 16'h2B05, 16'h280E, 
    16'h2526, 16'h224F, 16'h1F8B, 16'h1CDA, 16'h1A40, 16'h17BE, 16'h1555, 16'h1306, 
    16'h10D4, 16'h0EBF, 16'h0CC9, 16'h0AF3, 16'h093E, 16'h07AC, 16'h063D, 16'h04F2, 
    16'h03CC, 16'h02CC, 16'h01F2, 16'h013F, 16'h00B4, 16'h0050, 16'h0014, 16'h0000
};
localparam [15:0] HANN_256 [0:255] = '{
    16'h0000, 16'h0004, 16'h0013, 16'h002C, 16'h004F, 16'h007C, 16'h00B2, 16'h00F3, 
    16'h013D, 16'h0191, 16'h01EE, 16'h0256, 16'h02C6, 16'h0341, 16'h03C5, 16'h0452, 
    16'h04E8, 16'h0588, 16'h0631, 16'h06E2, 16'h079D, 16'h0860, 16'h092C, 16'h0A01, 
    16'h0ADE, 16'h0BC3, 16'h0CB0, 16'h0DA5, 16'h0EA2, 16'h0FA7, 16'h10B3, 16'h11C7, 
    16'h12E2, 16'h1404, 16'h152C, 16'h165C, 16'h1791, 16'h18CD, 16'h1A10, 16'h1B58, 
    16'h1CA5, 16'h1DF9, 16'h1F51, 16'h20AF, 16'h2211, 16'h2378, 16'h24E4, 16'h2654, 
    16'h27C7, 16'h293F, 16'h2ABA, 16'h2C38, 16'h2DBA, 16'h2F3E, 16'h30C5, 16'h324E, 
    16'h33D9, 16'h3567, 16'h36F6, 16'h3886, 16'h3A17, 16'h3BAA, 16'h3D3D, 16'h3ED0, 
    16'h4064, 16'h41F8, 16'h438B, 16'h451E, 16'h46B0, 16'h4840, 16'h49D0, 16'h4B5E, 
    16'h4CEB, 16'h4E75, 16'h4FFD, 16'h5183, 16'h5305, 16'h5485, 16'h5602, 16'h577B, 
    16'h58F1, 16'h5A63, 16'h5BD1, 16'h5D3A, 16'h5E9F, 16'h5FFF, 16'h615A, 16'h62B0, 
    16'h6400, 16'h654B, 16'h6690, 16'h67CF, 16'h6908, 16'h6A3B, 16'h6B67, 16'h6C8C, 
    16'h6DAA, 16'h6EC2, 16'h6FD2, 16'h70DA, 16'h71DB, 16'h72D4, 16'h73C6, 16'h74AF, 
    16'h7590, 16'h7669, 16'h7739, 16'h7800, 16'h78BF, 16'h7976, 16'h7A23, 16'h7AC7, 
    16'h7B62, 16'h7BF4, 16'h7C7C, 16'h7CFC, 16'h7D71, 16'h7DDD, 16'h7E40, 16'h7E98, 
    16'h7EE8, 16'h7F2D, 16'h7F68, 16'h7F9A, 16'h7FC2, 16'h7FDF, 16'h7FF3, 16'h7FFD, 
    16'h7FFD, 16'h7FF3, 16'h7FDF, 16'h7FC2, 16'h7F9A, 16'h7F68, 16'h7F2D, 16'h7EE8, 
    16'h7E98, 16'h7E40, 16'h7DDD, 16'h7D71, 16'h7CFC, 16'h7C7C, 16'h7BF4, 16'h7B62, 
    16'h7AC7, 16'h7A23, 16'h7976, 16'h78BF, 16'h7800, 16'h7739, 16'h7669, 16'h7590, 
    16'h74AF, 16'h73C6, 16'h72D4, 16'h71DB, 16'h70DA, 16'h6FD2, 16'h6EC2, 16'h6DAA, 
    16'h6C8C, 16'h6B67, 16'h6A3B, 16'h6908, 16'h67CF, 16'h6690, 16'h654B, 16'h6400, 
    16'h62B0, 16'h615A, 16'h5FFF, 16'h5E9F, 16'h5D3A, 16'h5BD1, 16'h5A63, 16'h58F1, 
    16'h577B, 16'h5602, 16'h5485, 16'h5305, 16'h5183, 16'h4FFD, 16'h4E75, 16'h4CEB, 
    16'h4B5E, 16'h49D0, 16'h4840, 16'h46B0, 16'h451E, 16'h438B, 16'h41F8, 16'h4064, 
    16'h3ED0, 16'h3D3D, 16'h3BAA, 16'h3A17, 16'h3886, 16'h36F6, 16'h3567, 16'h33D9, 
    16'h324E, 16'h30C5, 16'h2F3E, 16'h2DBA, 16'h2C38, 16'h2ABA, 16'h293F, 16'h27C7, 
    16'h2654, 16'h24E4, 16'h2378, 16'h2211, 16'h20AF, 16'h1F51, 16'h1DF9, 16'h1CA5, 
    16'h1B58, 16'h1A10, 16'h18CD, 16'h1791, 16'h165C, 16'h152C, 16'h1404, 16'h12E2, 
    16'h11C7, 16'h10B3, 16'h0FA7, 16'h0EA2, 16'h0DA5, 16'h0CB0, 16'h0BC3, 16'h0ADE, 
    16'h0A01, 16'h092C, 16'h0860, 16'h079D, 16'h06E2, 16'h0631, 16'h0588, 16'h04E8, 
    16'h0452, 16'h03C5, 16'h0341, 16'h02C6, 16'h0256, 16'h01EE, 16'h0191, 16'h013D, 
    16'h00F3, 16'h00B2, 16'h007C, 16'h004F, 16'h002C, 16'h0013, 16'h0004, 16'h0000
};
// 512点汉宁窗系数 (Q1.15格式)
localparam [15:0] HANN_512 [0:511] = '{
    16'h0000,16'h0001,16'h0004,16'h000B,16'h0013,16'h001E,16'h002C,16'h003C,16'h004F,16'h0064,16'h007B,16'h0095,16'h00B2,16'h00D0,16'h00F2,16'h0115,16'h013C,16'h0164,16'h018F,16'h01BD,16'h01EC,16'h021F,16'h0253,16'h028A,16'h02C4,16'h02FF,16'h033E,16'h037E,16'h03C1,16'h0406,16'h044E,16'h0497,16'h04E3,16'h0532,16'h0582,16'h05D5,16'h062B,16'h0682,16'h06DC,16'h0737,16'h0795,16'h07F6,16'h0858,16'h08BD,16'h0923,16'h098C,16'h09F7,16'h0A64,16'h0AD3,16'h0B44,16'h0BB7,16'h0C2D,16'h0CA4,16'h0D1D,16'h0D98,16'h0E15,16'h0E94,16'h0F15,16'h0F98,16'h101D,16'h10A3,16'h112C,16'h11B6,16'h1242,16'h12D0,16'h135F,16'h13F1,16'h1484,16'h1518,16'h15AF,16'h1647,16'h16E0,16'h177B,16'h1818,16'h18B6,16'h1956,16'h19F7,16'h1A9A,16'h1B3E,16'h1BE4,16'h1C8B,16'h1D33,16'h1DDD,16'h1E88,16'h1F35,16'h1FE2,16'h2091,16'h2141,16'h21F2,16'h22A5,16'h2358,16'h240D,16'h24C3,16'h257A,16'h2632,16'h26EA,16'h27A4,16'h285F,16'h291B,16'h29D7,16'h2A95,16'h2B53,16'h2C12,16'h2CD2,16'h2D92,16'h2E54,16'h2F16,16'h2FD8,16'h309B,16'h315F,16'h3224,16'h32E9,16'h33AE,16'h3474,16'h353A,16'h3601,16'h36C8,16'h3790,16'h3858,16'h3920,16'h39E8,16'h3AB1,16'h3B7A,16'h3C43,16'h3D0C,16'h3DD5,16'h3E9E,16'h3F68,16'h4031,16'h40FB,16'h41C4,16'h428E,16'h4357,16'h4420,16'h44E9,16'h45B2,16'h467A,16'h4742,16'h480A,16'h48D2,16'h4999,16'h4A60,16'h4B27,16'h4BED,16'h4CB3,16'h4D78,16'h4E3D,16'h4F01,16'h4FC4,16'h5087,16'h514A,16'h520B,16'h52CC,16'h538C,16'h544C,16'h550A,16'h55C8,16'h5685,16'h5741,16'h57FD,16'h58B7,16'h5970,16'h5A28,16'h5AE0,16'h5B96,16'h5C4B,16'h5CFF,16'h5DB2,16'h5E64,16'h5F15,16'h5FC5,16'h6073,16'h6120,16'h61CB,16'h6276,16'h631F,16'h63C7,16'h646D,16'h6512,16'h65B5,16'h6657,16'h66F8,16'h6797,16'h6835,16'h68D0,16'h696B,16'h6A04,16'h6A9B,16'h6B30,16'h6BC4,16'h6C56,16'h6CE7,16'h6D75,16'h6E02,16'h6E8D,16'h6F17,16'h6F9E,16'h7024,16'h70A7,16'h7129,16'h71A9,16'h7227,16'h72A4,16'h731E,16'h7396,16'h740C,16'h7480,16'h74F3,16'h7563,16'h75D1,16'h763D,16'h76A7,16'h770E,16'h7774,16'h77D7,16'h7839,16'h7898,16'h78F5,16'h7950,16'h79A8,16'h79FE,16'h7A52,16'h7AA4,16'h7AF4,16'h7B41,16'h7B8C,16'h7BD4,16'h7C1B,16'h7C5F,16'h7CA0,16'h7CE0,16'h7D1D,16'h7D57,16'h7D90,16'h7DC5,16'h7DF9,16'h7E2A,16'h7E58,16'h7E85,16'h7EAE,16'h7ED6,16'h7EFB,16'h7F1D,16'h7F3D,16'h7F5B,16'h7F76,16'h7F8F,16'h7FA5,16'h7FB9,16'h7FCA,16'h7FD9,16'h7FE5,16'h7FEF,16'h7FF7,16'h7FFC,16'h7FFE,16'h7FFE,16'h7FFC,16'h7FF7,16'h7FEF,16'h7FE5,16'h7FD9,16'h7FCA,16'h7FB9,16'h7FA5,16'h7F8F,16'h7F76,16'h7F5B,16'h7F3D,16'h7F1D,16'h7EFB,16'h7ED6,16'h7EAE,16'h7E85,16'h7E58,16'h7E2A,16'h7DF9,16'h7DC5,16'h7D90,16'h7D57,16'h7D1D,16'h7CE0,16'h7CA0,16'h7C5F,16'h7C1B,16'h7BD4,16'h7B8C,16'h7B41,16'h7AF4,16'h7AA4,16'h7A52,16'h79FE,16'h79A8,16'h7950,16'h78F5,16'h7898,16'h7839,16'h77D7,16'h7774,16'h770E,16'h76A7,16'h763D,16'h75D1,16'h7563,16'h74F3,16'h7480,16'h740C,16'h7396,16'h731E,16'h72A4,16'h7227,16'h71A9,16'h7129,16'h70A7,16'h7024,16'h6F9E,16'h6F17,16'h6E8D,16'h6E02,16'h6D75,16'h6CE7,16'h6C56,16'h6BC4,16'h6B30,16'h6A9B,16'h6A04,16'h696B,16'h68D0,16'h6835,16'h6797,16'h66F8,16'h6657,16'h65B5,16'h6512,16'h646D,16'h63C7,16'h631F,16'h6276,16'h61CB,16'h6120,16'h6073,16'h5FC5,16'h5F15,16'h5E64,16'h5DB2,16'h5CFF,16'h5C4B,16'h5B96,16'h5AE0,16'h5A28,16'h5970,16'h58B7,16'h57FD,16'h5741,16'h5685,16'h55C8,16'h550A,16'h544C,16'h538C,16'h52CC,16'h520B,16'h514A,16'h5087,16'h4FC4,16'h4F01,16'h4E3D,16'h4D78,16'h4CB3,16'h4BED,16'h4B27,16'h4A60,16'h4999,16'h48D2,16'h480A,16'h4742,16'h467A,16'h45B2,16'h44E9,16'h4420,16'h4357,16'h428E,16'h41C4,16'h40FB,16'h4031,16'h3F68,16'h3E9E,16'h3DD5,16'h3D0C,16'h3C43,16'h3B7A,16'h3AB1,16'h39E8,16'h3920,16'h3858,16'h3790,16'h36C8,16'h3601,16'h353A,16'h3474,16'h33AE,16'h32E9,16'h3224,16'h315F,16'h309B,16'h2FD8,16'h2F16,16'h2E54,16'h2D92,16'h2CD2,16'h2C12,16'h2B53,16'h2A95,16'h29D7,16'h291B,16'h285F,16'h27A4,16'h26EA,16'h2632,16'h257A,16'h24C3,16'h240D,16'h2358,16'h22A5,16'h21F2,16'h2141,16'h2091,16'h1FE2,16'h1F35,16'h1E88,16'h1DDD,16'h1D33,16'h1C8B,16'h1BE4,16'h1B3E,16'h1A9A,16'h19F7,16'h1956,16'h18B6,16'h1818,16'h177B,16'h16E0,16'h1647,16'h15AF,16'h1518,16'h1484,16'h13F1,16'h135F,16'h12D0,16'h1242,16'h11B6,16'h112C,16'h10A3,16'h101D,16'h0F98,16'h0F15,16'h0E94,16'h0E15,16'h0D98,16'h0D1D,16'h0CA4,16'h0C2D,16'h0BB7,16'h0B44,16'h0AD3,16'h0A64,16'h09F7,16'h098C,16'h0923,16'h08BD,16'h0858,16'h07F6,16'h0795,16'h0737,16'h06DC,16'h0682,16'h062B,16'h05D5,16'h0582,16'h0532,16'h04E3,16'h0497,16'h044E,16'h0406,16'h03C1,16'h037E,16'h033E,16'h02FF,16'h02C4,16'h028A,16'h0253,16'h021F,16'h01EC,16'h01BD,16'h018F,16'h0164,16'h013C,16'h0115,16'h00F2,16'h00D0,16'h00B2,16'h0095,16'h007B,16'h0064,16'h004F,16'h003C,16'h002C,16'h001E,16'h0013,16'h000B,16'h0004,16'h0001,16'h0000
};

endpackage

`endif // HANN_WINDOW_COEFF_SV